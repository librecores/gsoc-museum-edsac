module ccu_4
  (output reg ep3,
   output reg g6_pos,

   input wire c1,
   input wire ev_d0,
   input wire g8,
   input wire odd_d0,
   input wire r2);

   // Body

endmodule // ccu_4
