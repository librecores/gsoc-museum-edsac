module order_tank
  (output reg gated_order,
   output reg ungated_order,

   input wire clk,
   input wire cu_gate_pos,
   input wire eng_mode_neg,
   input wire eng_order,
   input wire epsep,
   input wire g12,
   input wire mob,
   input wire clr_order,
   input wire starter_neg);

   // Contains one half cycle delay line.

   // Body

endmodule // order_tank
