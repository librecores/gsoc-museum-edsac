module coincidence
  (output reg cu_gate_pos,
   output reg cu_gate_neg,
   output reg order_sct,
   output reg r_pulse,

   input wire cntr,
   input wire d0,
   input wire d2,
   input wire d7,
   input wire d18,
   input wire d20,
   input wire d25,
   input wire f1_neg,
   input wire order,
   input wire s1,
   input wire sct);

   // Body

endmodule // coincidence
