module order_decoder2_1
  (output reg op_erase,
   output reg op_i,
   output reg op_j,
   output reg op_k,
   output reg op_o,
   output reg op_pi,
   output reg op_s,
   output reg op_z,

   input wire f13_pos,
   input wire f13_neg,
   input wire f14_pos,
   input wire f14_neg,
   input wire f15_pos,
   input wire f15_neg,
   input wire o_dy_1);

   // One order_decoder2 to be instantiated.

endmodule // order_decoder2_1
