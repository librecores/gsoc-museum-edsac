module ccu_8
  (output reg ep1,
   output reg g4_pos,
   output reg g4_neg,
   output reg ones2,

   input wire seventy_d35,
   input wire c11,
   input wire c14,
   input wire da,
   input wire ds_r,
   input wire dy,
   input wire ep_done,
   input wire ev_d0,
   input wire odd_d35,
   input wire g5,
   input wire reset_shift_ff);

   // Body

endmodule // ccu_8
