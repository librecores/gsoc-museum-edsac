module acc_shift_ii
  (output reg adder_a,

   input wire clk,
   input wire acc1,
   input wire x1,
   input wire x2,
   input wire x3,
   input wire x4);

   // Body

endmodule // acc_shift_ii
