/* Module for Starter Unit/Initial Orders Loader.
 */

module starter (
  output wire boot_valid,
  output wire ep9,
  output wire reset_cntr_neg,
  output wire reset_sct_neg,
  output wire mob_starter,
  output wire sep2,
  output wire starter,
  output wire starter_neg,
  output wire stop_one_d,

  input wire  initial_orders, // Serial input of initial orders.
  input wire  s2,
  input wire  start,
  input wire  d17,
  input wire  d18,
  input wire  d19,
  input wire  d20,
  input wire  d21,
  input wire  d22,
  input wire  d23,
  input wire  d24,
  input wire  d25,
  input wire  d26,
  input wire  d27,
  input wire  d28,
  input wire  d29,
  input wire  d30,
  input wire  d31,
  input wire  d32,
  input wire  d33,
  input wire  d34,
  input wire  d35
  );

endmodule
