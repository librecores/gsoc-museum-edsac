/* Module for Engineers Control Panel.
 */

module engineer_control_panel (
  output wire eng_mode_neg,
  output wire eng_order,
  output wire order_clr,

  input wire  d0,
  input wire  d18,
  input wire  d19,
  input wire  d20,
  input wire  d21,
  input wire  d22,
  input wire  d23,
  input wire  d24,
  input wire  d25,
  input wire  d26,
  input wire  d27,
  input wire  d28,
  input wire  d29,
  input wire  d30,
  input wire  d31,
  input wire  d32,
  input wire  d33,
  input wire  d34,
  input wire  d35,
  input wire  o1_t_btn,
  input wire  o2_t_btn,
  input wire  o3_t_btn,
  input wire  o4_t_btn,
  input wire  o5_t_btn,
  input wire  o6_t_btn,
  input wire  o7_t_btn,
  input wire  o8_t_btn,
  input wire  o9_t_btn,
  input wire  o10_t_btn,
  input wire  o11_t_btn,
  input wire  o12_t_btn,
  input wire  o13_t_btn,
  input wire  o14_t_btn,
  input wire  o15_t_btn,
  input wire  o16_t_btn,
  input wire  o17_t_btn,
  input wire  eng_mode_t_btn
  );

endmodule
