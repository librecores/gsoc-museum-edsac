module ccu_3
  (output reg ep2,
   output reg g5,
   output reg reset_shift_ff,

   input wire zero_d0,
   input wire c6,
   input wire dy,
   input wire ev_d0,
   input wire ev_d1,
   input wire ungated_order);

   // Body

endmodule // ccu_3
