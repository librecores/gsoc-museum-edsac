module memory_f1_up_0
  (output reg monitor1,
   output reg f1_up_mob_t0,

   input wire f1_clk,
   input wire f1_mib,
   input wire f1_up_t0_clr,
   input wire f1_up_t0_in,
   input wire f1_up_t0_out);

   // Atomic dleay_line module to be instantiated here 
   // with 1.152ms delay for circulation of 16 full 
   // words or 32 short words (instructions).

   // Body

endmodule // memory_f1_up_0
