module transfer (
  output wire mib,
  output wire mob,

  input wire  clk,
  input wire  f1_pos,
  input wire  f2_pos,
  input wire  mob_asu1,
  input wire  mob_tape,
  input wire  mob_starter,
  input wire  mob_printer,
  input wire  f1_mob,
  input wire  f2_mob,
  input wire  r1_mob,
  input wire  r2_mob
  );

  // Body

endmodule // transfer
