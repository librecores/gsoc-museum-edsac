module counter
  (output reg cntr,

   input wire clk,
   input wire d1,
   input wire d19,
   input wire reset_cntr);

   // One half adder to be instantiated 
   // along with half cycle delay.

   // Body

endmodule // counter
