/* Top Level L0 EDSAC module.
 */

module edsac (
  input wire clk,
  // Push buttons.
  input wire resume_btn,
  input wire single_ep_btn,
  input wire start_btn,
  input wire stop_btn,
  input wire extended_btn,
  // Toggle buttons.
  input wire o1_t_btn,
  input wire o2_t_btn,
  input wire o3_t_btn,
  input wire o4_t_btn,
  input wire o5_t_btn,
  input wire o6_t_btn,
  input wire o7_t_btn,
  input wire o8_t_btn,
  input wire o9_t_btn,
  input wire o10_t_btn,
  input wire o11_t_btn,
  input wire o12_t_btn,
  input wire o13_t_btn,
  input wire o14_t_btn,
  input wire o15_t_btn,
  input wire o16_t_btn,
  input wire o17_t_btn,
  input wire eng_mode_t_btn
  );

  wire        f1_down_mob_t0;
  wire        f1_up_mob_t0;
  wire        f1_down_mob_t1;
  wire        f1_up_mob_t1;
  wire        f1_down_mob_t2;
  wire        f1_up_mob_t2;
  wire        f1_down_mob_t3;
  wire        f1_up_mob_t3;
  wire        f2_down_mob_t0;
  wire        f2_up_mob_t0;
  wire        f2_down_mob_t1;
  wire        f2_up_mob_t1;
  wire        f2_down_mob_t2;
  wire        f2_up_mob_t2;
  wire        f2_down_mob_t3;
  wire        f2_up_mob_t3;
  wire        r1_down_mob_t0;
  wire        r1_up_mob_t0;
  wire        r1_down_mob_t1;
  wire        r1_up_mob_t1;
  wire        r1_down_mob_t2;
  wire        r1_up_mob_t2;
  wire        r1_down_mob_t3;
  wire        r1_up_mob_t3;
  wire        r2_down_mob_t0;
  wire        r2_up_mob_t0;
  wire        r2_down_mob_t1;
  wire        r2_up_mob_t1;
  wire        r2_down_mob_t2;
  wire        r2_up_mob_t2;
  wire        r2_down_mob_t3;
  wire        r2_up_mob_t3;
  wire        f1_mib;
  wire        f2_mib;
  wire        r1_mib;
  wire        r2_mib;
  wire        f1_down_t0_clr;
  wire        f1_up_t0_clr;
  wire        f1_down_t1_clr;
  wire        f1_up_t1_clr;
  wire        f1_down_t2_clr;
  wire        f1_up_t2_clr;
  wire        f1_down_t3_clr;
  wire        f1_up_t3_clr;
  wire        f2_down_t0_clr;
  wire        f2_up_t0_clr;
  wire        f2_down_t1_clr;
  wire        f2_up_t1_clr;
  wire        f2_down_t2_clr;
  wire        f2_up_t2_clr;
  wire        f2_down_t3_clr;
  wire        f2_up_t3_clr;
  wire        r1_down_t0_clr;
  wire        r1_up_t0_clr;
  wire        r1_down_t1_clr;
  wire        r1_up_t1_clr;
  wire        r1_down_t2_clr;
  wire        r1_up_t2_clr;
  wire        r1_down_t3_clr;
  wire        r1_up_t3_clr;
  wire        r2_down_t0_clr;
  wire        r2_up_t0_clr;
  wire        r2_down_t1_clr;
  wire        r2_up_t1_clr;
  wire        r2_down_t2_clr;
  wire        r2_up_t2_clr;
  wire        r2_down_t3_clr;
  wire        r2_up_t3_clr;
  wire        f1_up_t0_in;
  wire        f1_up_t1_in;
  wire        f1_up_t2_in;
  wire        f1_up_t3_in;
  wire        f1_down_t0_in;
  wire        f1_down_t1_in;
  wire        f1_down_t2_in;
  wire        f1_down_t3_in;
  wire        f1_up_t0_out;
  wire        f1_up_t1_out;
  wire        f1_up_t2_out;
  wire        f1_up_t3_out;
  wire        f1_down_t0_out;
  wire        f1_down_t1_out;
  wire        f1_down_t2_out;
  wire        f1_down_t3_out;
  wire        f2_up_t0_in;
  wire        f2_up_t1_in;
  wire        f2_up_t2_in;
  wire        f2_up_t3_in;
  wire        f2_down_t0_in;
  wire        f2_down_t1_in;
  wire        f2_down_t2_in;
  wire        f2_down_t3_in;
  wire        f2_up_t0_out;
  wire        f2_up_t1_out;
  wire        f2_up_t2_out;
  wire        f2_up_t3_out;
  wire        f2_down_t0_out;
  wire        f2_down_t1_out;
  wire        f2_down_t2_out;
  wire        f2_down_t3_out;
  wire        r1_up_t0_in;
  wire        r1_up_t1_in;
  wire        r1_up_t2_in;
  wire        r1_up_t3_in;
  wire        r1_down_t0_in;
  wire        r1_down_t1_in;
  wire        r1_down_t2_in;
  wire        r1_down_t3_in;
  wire        r1_up_t0_out;
  wire        r1_up_t1_out;
  wire        r1_up_t2_out;
  wire        r1_up_t3_out;
  wire        r1_down_t0_out;
  wire        r1_down_t1_out;
  wire        r1_down_t2_out;
  wire        r1_down_t3_out;
  wire        r2_up_t0_in;
  wire        r2_up_t1_in;
  wire        r2_up_t2_in;
  wire        r2_up_t3_in;
  wire        r2_down_t0_in;
  wire        r2_down_t1_in;
  wire        r2_down_t2_in;
  wire        r2_down_t3_in;
  wire        r2_up_t0_out;
  wire        r2_up_t1_out;
  wire        r2_up_t2_out;
  wire        r2_up_t3_out;
  wire        r2_down_t0_out;
  wire        r2_down_t1_out;
  wire        r2_down_t2_out;
  wire        r2_down_t3_out;
  wire [35:0] d;
  wire        mcand_in;
  wire        da_n;
  wire        dx_m;
  wire        ep4;
  wire        ds_r;
  wire        dv_d;
  wire        mob;
  wire        mib;
  wire        c1;
  wire        c2;
  wire        c3;
  wire        c4;
  wire        c7;
  wire        c8;
  wire        c9;
  wire        c10;
  wire        c18;
  wire        c19;
  wire        c21;
  wire        c25;
  wire        g12;
  wire        g13;
  wire        r2;
  wire        g2_pos;
  wire        g2_neg;
  wire        dx;
  wire        g1_pos;
  wire        g1_neg;
  wire        g3_pos;
  wire        g4_pos;
  wire        g4_neg;
  wire        g5;
  wire        g6_pos;
  wire        g9_neg;
  wire        g10_neg;
  wire        g11_neg;
  wire        da_m;
  wire        ccu_ones;
  wire        ev_d1_dz;
  wire        ds;
  wire        dv;
  wire        jump_uc;
  wire        f1_neg;
  wire        s2;
  wire        ep9;
  wire        reset_cntr_neg;
  wire        starter;
  wire        starter_neg;
  wire        reset_sct_neg;
  wire        ev_d1;
  wire        ep_done;
  wire        ep10;
  wire        ep8;
  wire        stop_one_a;
  wire        stop_one_c;
  wire        c16;
  wire        mob_asu1;
  wire        mob_tape;
  wire        mob_starter;
  wire        mob_printer;
  wire        epsep;
  wire        ep11;
  wire        extended_pos;
  wire        extended_neg;
  wire        single_ep;
  wire        start;
  wire        stop_neg;
  wire        c22;
  wire        ep;
  wire        sep2;

  computer computer (
    .mcand_in (mcand_in),
    .da_n     (da_n),
    .dx_m     (dx_m),
    .ep4      (ep4),
    .ds_r     (ds_r),
    .dv_d     (dv_d),
    .mob      (mob),
    .mib      (mib),
    .clk      (clk),
    .d0       (d[0]),
    .d17      (d[17]),
    .d35      (d[35]),
    .c1       (c1),
    .c2       (c2),
    .c3       (c3),
    .c4       (c4),
    .c7       (c7),
    .c8       (c8),
    .c9       (c9),
    .c10      (c10),
    .c18      (c18),
    .c19      (c19),
    .c21      (c21),
    .c25      (c25),
    .g12      (g12),
    .g13      (g13),
    .r2       (r2),
    .g2_pos   (g2_pos),
    .g2_neg   (g2_neg),
    .dx       (dx),
    .g1_pos   (g1_pos),
    .g1_neg   (g1_neg),
    .g3_pos   (g3_pos),
    .g4_pos   (g4_pos),
    .g4_neg   (g4_neg),
    .g5       (g5),
    .g6_pos   (g6_pos),
    .g9_neg   (g9_neg),
    .g10_neg  (g10_neg),
    .g11_neg  (g11_neg),
    .da_m     (da_m),
    .ccu_ones (ccu_ones),
    .ev_d1_dz (ev_d1_dz),
    .ds       (ds),
    .dv       (dv),
    .jump_uc  (jump_uc),
    .f1_neg   (f1_neg)
    );

  control_section control_section (
    .s2             (s2),
    .ep9            (ep9),
    .reset_cntr_neg (reset_cntr_neg),
    .starter        (starter),
    .starter_neg    (starter_neg),
    .reset_sct_neg  (reset_sct_neg),
    .g1_pos         (g1_pos),
    .g1_neg         (g1_neg),
    .ev_d1_dz       (ev_d1_dz),
    .ev_d1          (ev_d1),
    .da_m           (da_m),
    .ds             (ds),
    .g5             (g5),
    .g6_pos         (g6_pos),
    .ccu_ones       (ccu_ones),
    .g2_pos         (g2_pos),
    .g2_neg         (g2_neg),
    .g3_pos         (g3_pos),
    .g4_pos         (g4_pos),
    .g4_neg         (g4_neg),
    .g9_neg         (g9_neg),
    .g10_neg        (g10_neg),
    .g11_neg        (g11_neg),
    .dv             (dv),
    .jump_uc        (jump_uc),
    .r2             (r2),
    .g12            (g12),
    .g13            (g13),
    .f1_neg         (f1_neg),
    .mib            (mib),
    .mcand_in       (mcand_in),
    .da_n           (da_n),
    .ds_r           (ds_r),
    .ep4            (ep4),
    .dx_m           (dx_m),
    .dv_d           (dv_d),
    .dx             (dx),
    .d0             (d[0]),
    .d1             (d[1]),
    .d2             (d[2]),
    .d7             (d[7]),
    .d18            (d[18]),
    .d19            (d[19]),
    .d20            (d[20]),
    .d21            (d[21]),
    .d22            (d[22]),
    .d23            (d[23]),
    .d24            (d[24]),
    .d25            (d[25]),
    .d26            (d[26]),
    .d27            (d[27]),
    .d28            (d[28]),
    .d29            (d[29]),
    .d31            (d[31]),
    .d32            (d[32]),
    .d33            (d[33]),
    .d34            (d[34]),
    .d35            (d[35]),
    .ep_done        (ep_done),
    .ep10           (ep10),
    .ep8            (ep8),
    .stop_one_a     (stop_one_a),
    .stop_one_c     (stop_one_c),
    .c1             (c1),
    .c2             (c2),
    .c3             (c3),
    .c4             (c4),
    .c7             (c7),
    .c8             (c8),
    .c9             (c9),
    .c10            (c10),
    .c16            (c16),
    .c18            (c18),
    .c19            (c19),
    .c21            (c21),
    .c25            (c25),
    .f1_down_t0_clr (f1_down_t0_clr),
    .f1_up_t0_clr   (f1_up_t0_clr),
    .f1_down_t1_clr (f1_down_t1_clr),
    .f1_up_t1_clr   (f1_up_t1_clr),
    .f1_down_t2_clr (f1_down_t2_clr),
    .f1_up_t2_clr   (f1_up_t2_clr),
    .f1_down_t3_clr (f1_down_t3_clr),
    .f1_up_t3_clr   (f1_up_t3_clr),
    .f2_down_t0_clr (f2_down_t0_clr),
    .f2_up_t0_clr   (f2_up_t0_clr),
    .f2_down_t1_clr (f2_down_t1_clr),
    .f2_up_t1_clr   (f2_up_t1_clr),
    .f2_down_t2_clr (f2_down_t2_clr),
    .f2_up_t2_clr   (f2_up_t2_clr),
    .f2_down_t3_clr (f2_down_t3_clr),
    .f2_up_t3_clr   (f2_up_t3_clr),
    .r1_down_t0_clr (r1_down_t0_clr),
    .r1_up_t0_clr   (r1_up_t0_clr),
    .r1_down_t1_clr (r1_down_t1_clr),
    .r1_up_t1_clr   (r1_up_t1_clr),
    .r1_down_t2_clr (r1_down_t2_clr),
    .r1_up_t2_clr   (r1_up_t2_clr),
    .r1_down_t3_clr (r1_down_t3_clr),
    .r1_up_t3_clr   (r1_up_t3_clr),
    .r2_down_t0_clr (r2_down_t0_clr),
    .r2_up_t0_clr   (r2_up_t0_clr),
    .r2_down_t1_clr (r2_down_t1_clr),
    .r2_up_t1_clr   (r2_up_t1_clr),
    .r2_down_t2_clr (r2_down_t2_clr),
    .r2_up_t2_clr   (r2_up_t2_clr),
    .r2_down_t3_clr (r2_down_t3_clr),
    .r2_up_t3_clr   (r2_up_t3_clr),
    .f1_mib         (f1_mib),
    .f2_mib         (f2_mib),
    .r1_mib         (r1_mib),
    .r2_mib         (r2_mib),
    .f1_up_t0_in    (f1_up_t0_in),
    .f1_up_t1_in    (f1_up_t1_in),
    .f1_up_t2_in    (f1_up_t2_in),
    .f1_up_t3_in    (f1_up_t3_in),
    .f1_down_t0_in  (f1_down_t0_in),
    .f1_down_t1_in  (f1_down_t1_in),
    .f1_down_t2_in  (f1_down_t2_in),
    .f1_down_t3_in  (f1_down_t3_in),
    .f1_up_t0_out   (f1_up_t0_out),
    .f1_up_t1_out   (f1_up_t1_out),
    .f1_up_t2_out   (f1_up_t2_out),
    .f1_up_t3_out   (f1_up_t3_out),
    .f1_down_t0_out (f1_down_t0_out),
    .f1_down_t1_out (f1_down_t1_out),
    .f1_down_t2_out (f1_down_t2_out),
    .f1_down_t3_out (f1_down_t3_out),
    .f2_up_t0_in    (f2_up_t0_in),
    .f2_up_t1_in    (f2_up_t1_in),
    .f2_up_t2_in    (f2_up_t2_in),
    .f2_up_t3_in    (f2_up_t3_in),
    .f2_down_t0_in  (f2_down_t0_in),
    .f2_down_t1_in  (f2_down_t1_in),
    .f2_down_t2_in  (f2_down_t2_in),
    .f2_down_t3_in  (f2_down_t3_in),
    .f2_up_t0_out   (f2_up_t0_out),
    .f2_up_t1_out   (f2_up_t1_out),
    .f2_up_t2_out   (f2_up_t2_out),
    .f2_up_t3_out   (f2_up_t3_out),
    .f2_down_t0_out (f2_down_t0_out),
    .f2_down_t1_out (f2_down_t1_out),
    .f2_down_t2_out (f2_down_t2_out),
    .f2_down_t3_out (f2_down_t3_out),
    .r1_up_t0_in    (r1_up_t0_in),
    .r1_up_t1_in    (r1_up_t1_in),
    .r1_up_t2_in    (r1_up_t2_in),
    .r1_up_t3_in    (r1_up_t3_in),
    .r1_down_t0_in  (r1_down_t0_in),
    .r1_down_t1_in  (r1_down_t1_in),
    .r1_down_t2_in  (r1_down_t2_in),
    .r1_down_t3_in  (r1_down_t3_in),
    .r1_up_t0_out   (r1_up_t0_out),
    .r1_up_t1_out   (r1_up_t1_out),
    .r1_up_t2_out   (r1_up_t2_out),
    .r1_up_t3_out   (r1_up_t3_out),
    .r1_down_t0_out (r1_down_t0_out),
    .r1_down_t1_out (r1_down_t1_out),
    .r1_down_t2_out (r1_down_t2_out),
    .r1_down_t3_out (r1_down_t3_out),
    .r2_up_t0_in    (r2_up_t0_in),
    .r2_up_t1_in    (r2_up_t1_in),
    .r2_up_t2_in    (r2_up_t2_in),
    .r2_up_t3_in    (r2_up_t3_in),
    .r2_down_t0_in  (r2_down_t0_in),
    .r2_down_t1_in  (r2_down_t1_in),
    .r2_down_t2_in  (r2_down_t2_in),
    .r2_down_t3_in  (r2_down_t3_in),
    .r2_up_t0_out   (r2_up_t0_out),
    .r2_up_t1_out   (r2_up_t1_out),
    .r2_up_t2_out   (r2_up_t2_out),
    .r2_up_t3_out   (r2_up_t3_out),
    .r2_down_t0_out (r2_down_t0_out),
    .r2_down_t1_out (r2_down_t1_out),
    .r2_down_t2_out (r2_down_t2_out),
    .r2_down_t3_out (r2_down_t3_out),
    .f1_down_mob_t0 (f1_down_mob_t0),
    .f1_up_mob_t0   (f1_up_mob_t0),
    .f1_down_mob_t1 (f1_down_mob_t1),
    .f1_up_mob_t1   (f1_up_mob_t1),
    .f1_down_mob_t2 (f1_down_mob_t2),
    .f1_up_mob_t2   (f1_up_mob_t2),
    .f1_down_mob_t3 (f1_down_mob_t3),
    .f1_up_mob_t3   (f1_up_mob_t3),
    .f2_down_mob_t0 (f2_down_mob_t0),
    .f2_up_mob_t0   (f2_up_mob_t0),
    .f2_down_mob_t1 (f2_down_mob_t1),
    .f2_up_mob_t1   (f2_up_mob_t1),
    .f2_down_mob_t2 (f2_down_mob_t2),
    .f2_up_mob_t2   (f2_up_mob_t2),
    .f2_down_mob_t3 (f2_down_mob_t3),
    .f2_up_mob_t3   (f2_up_mob_t3),
    .r1_down_mob_t0 (r1_down_mob_t0),
    .r1_up_mob_t0   (r1_up_mob_t0),
    .r1_down_mob_t1 (r1_down_mob_t1),
    .r1_up_mob_t1   (r1_up_mob_t1),
    .r1_down_mob_t2 (r1_down_mob_t2),
    .r1_up_mob_t2   (r1_up_mob_t2),
    .r1_down_mob_t3 (r1_down_mob_t3),
    .r1_up_mob_t3   (r1_up_mob_t3),
    .r2_down_mob_t0 (r2_down_mob_t0),
    .r2_up_mob_t0   (r2_up_mob_t0),
    .r2_down_mob_t1 (r2_down_mob_t1),
    .r2_up_mob_t1   (r2_up_mob_t1),
    .r2_down_mob_t2 (r2_down_mob_t2),
    .r2_up_mob_t2   (r2_up_mob_t2),
    .r2_down_mob_t3 (r2_down_mob_t3),
    .r2_up_mob_t3   (r2_up_mob_t3),
    .mob_asu1       (mob_asu1),
    .mob_tape       (mob_tape),
    .mob_starter    (mob_starter),
    .mob_printer    (mob_printer),
    .o1_t_btn       (o1_t_btn),
    .o2_t_btn       (o2_t_btn),
    .o3_t_btn       (o3_t_btn),
    .o4_t_btn       (o4_t_btn),
    .o5_t_btn       (o5_t_btn),
    .o6_t_btn       (o6_t_btn),
    .o7_t_btn       (o7_t_btn),
    .o8_t_btn       (o8_t_btn),
    .o9_t_btn       (o9_t_btn),
    .o10_t_btn      (o10_t_btn),
    .o11_t_btn      (o11_t_btn),
    .o12_t_btn      (o12_t_btn),
    .o13_t_btn      (o13_t_btn),
    .o14_t_btn      (o14_t_btn),
    .o15_t_btn      (o15_t_btn),
    .o16_t_btn      (o16_t_btn),
    .o17_t_btn      (o17_t_btn),
    .eng_mode_t_btn (eng_mode_t_btn)
    );

  digit_pulse_generator digit_pulse_generator (
    .digit_pulse (d[35:0]),
    
    .clk (clk)
    );

  memory_top memory_top (
    // TODO: monitors are for displaying Tank contents and are not connected for now.
    .monitor1       (),
    .monitor2       (),
    .monitor3       (),
    .monitor4       (),
    .monitor5       (),
    .monitor6       (),
    .monitor7       (),
    .monitor8       (),
    .monitor9       (),
    .monitor10      (),
    .monitor11      (),
    .monitor12      (),
    .monitor13      (),
    .monitor14      (),
    .monitor15      (),
    .monitor16      (),
    .monitor17      (),
    .monitor18      (),
    .monitor19      (),
    .monitor20      (),
    .monitor21      (),
    .monitor22      (),
    .monitor23      (),
    .monitor24      (),
    .monitor25      (),
    .monitor26      (),
    .monitor27      (),
    .monitor28      (),
    .monitor29      (),
    .monitor30      (),
    .monitor31      (),
    .monitor32      (),
    .f1_down_mob_t0 (f1_down_mob_t0),
    .f1_up_mob_t0   (f1_up_mob_t0),
    .f1_down_mob_t1 (f1_down_mob_t1),
    .f1_up_mob_t1   (f1_up_mob_t1),
    .f1_down_mob_t2 (f1_down_mob_t2),
    .f1_up_mob_t2   (f1_up_mob_t2),
    .f1_down_mob_t3 (f1_down_mob_t3),
    .f1_up_mob_t3   (f1_up_mob_t3),
    .f2_down_mob_t0 (f2_down_mob_t0),
    .f2_up_mob_t0   (f2_up_mob_t0),
    .f2_down_mob_t1 (f2_down_mob_t1),
    .f2_up_mob_t1   (f2_up_mob_t1),
    .f2_down_mob_t2 (f2_down_mob_t2),
    .f2_up_mob_t2   (f2_up_mob_t2),
    .f2_down_mob_t3 (f2_down_mob_t3),
    .f2_up_mob_t3   (f2_up_mob_t3),
    .r1_down_mob_t0 (r1_down_mob_t0),
    .r1_up_mob_t0   (r1_up_mob_t0),
    .r1_down_mob_t1 (r1_down_mob_t1),
    .r1_up_mob_t1   (r1_up_mob_t1),
    .r1_down_mob_t2 (r1_down_mob_t2),
    .r1_up_mob_t2   (r1_up_mob_t2),
    .r1_down_mob_t3 (r1_down_mob_t3),
    .r1_up_mob_t3   (r1_up_mob_t3),
    .r2_down_mob_t0 (r2_down_mob_t0),
    .r2_up_mob_t0   (r2_up_mob_t0),
    .r2_down_mob_t1 (r2_down_mob_t1),
    .r2_up_mob_t1   (r2_up_mob_t1),
    .r2_down_mob_t2 (r2_down_mob_t2),
    .r2_up_mob_t2   (r2_up_mob_t2),
    .r2_down_mob_t3 (r2_down_mob_t3),
    .r2_up_mob_t3   (r2_up_mob_t3),

    .f1_mib         (f1_mib),
    .f2_mib         (f2_mib),
    .r1_mib         (r1_mib),
    .r2_mib         (r2_mib),
    .f1_down_t0_clr (f1_down_t0_clr),
    .f1_up_t0_clr   (f1_up_t0_clr),
    .f1_down_t1_clr (f1_down_t1_clr),
    .f1_up_t1_clr   (f1_up_t1_clr),
    .f1_down_t2_clr (f1_down_t2_clr),
    .f1_up_t2_clr   (f1_up_t2_clr),
    .f1_down_t3_clr (f1_down_t3_clr),
    .f1_up_t3_clr   (f1_up_t3_clr),
    .f2_down_t0_clr (f2_down_t0_clr),
    .f2_up_t0_clr   (f2_up_t0_clr),
    .f2_down_t1_clr (f2_down_t1_clr),
    .f2_up_t1_clr   (f2_up_t1_clr),
    .f2_down_t2_clr (f2_down_t2_clr),
    .f2_up_t2_clr   (f2_up_t2_clr),
    .f2_down_t3_clr (f2_down_t3_clr),
    .f2_up_t3_clr   (f2_up_t3_clr),
    .r1_down_t0_clr (r1_down_t0_clr),
    .r1_up_t0_clr   (r1_up_t0_clr),
    .r1_down_t1_clr (r1_down_t1_clr),
    .r1_up_t1_clr   (r1_up_t1_clr),
    .r1_down_t2_clr (r1_down_t2_clr),
    .r1_up_t2_clr   (r1_up_t2_clr),
    .r1_down_t3_clr (r1_down_t3_clr),
    .r1_up_t3_clr   (r1_up_t3_clr),
    .r2_down_t0_clr (r2_down_t0_clr),
    .r2_up_t0_clr   (r2_up_t0_clr),
    .r2_down_t1_clr (r2_down_t1_clr),
    .r2_up_t1_clr   (r2_up_t1_clr),
    .r2_down_t2_clr (r2_down_t2_clr),
    .r2_up_t2_clr   (r2_up_t2_clr),
    .r2_down_t3_clr (r2_down_t3_clr),
    .r2_up_t3_clr   (r2_up_t3_clr),
    .f1_up_t0_in    (f1_up_t0_in),
    .f1_up_t1_in    (f1_up_t1_in),
    .f1_up_t2_in    (f1_up_t2_in),
    .f1_up_t3_in    (f1_up_t3_in),
    .f1_down_t0_in  (f1_down_t0_in),
    .f1_down_t1_in  (f1_down_t1_in),
    .f1_down_t2_in  (f1_down_t2_in),
    .f1_down_t3_in  (f1_down_t3_in),
    .f1_up_t0_out   (f1_up_t0_out),
    .f1_up_t1_out   (f1_up_t1_out),
    .f1_up_t2_out   (f1_up_t2_out),
    .f1_up_t3_out   (f1_up_t3_out),
    .f1_down_t0_out (f1_down_t0_out),
    .f1_down_t1_out (f1_down_t1_out),
    .f1_down_t2_out (f1_down_t2_out),
    .f1_down_t3_out (f1_down_t3_out),
    .f2_up_t0_in    (f2_up_t0_in),
    .f2_up_t1_in    (f2_up_t1_in),
    .f2_up_t2_in    (f2_up_t2_in),
    .f2_up_t3_in    (f2_up_t3_in),
    .f2_down_t0_in  (f2_down_t0_in),
    .f2_down_t1_in  (f2_down_t1_in),
    .f2_down_t2_in  (f2_down_t2_in),
    .f2_down_t3_in  (f2_down_t3_in),
    .f2_up_t0_out   (f2_up_t0_out),
    .f2_up_t1_out   (f2_up_t1_out),
    .f2_up_t2_out   (f2_up_t2_out),
    .f2_up_t3_out   (f2_up_t3_out),
    .f2_down_t0_out (f2_down_t0_out),
    .f2_down_t1_out (f2_down_t1_out),
    .f2_down_t2_out (f2_down_t2_out),
    .f2_down_t3_out (f2_down_t3_out),
    .r1_up_t0_in    (r1_up_t0_in),
    .r1_up_t1_in    (r1_up_t1_in),
    .r1_up_t2_in    (r1_up_t2_in),
    .r1_up_t3_in    (r1_up_t3_in),
    .r1_down_t0_in  (r1_down_t0_in),
    .r1_down_t1_in  (r1_down_t1_in),
    .r1_down_t2_in  (r1_down_t2_in),
    .r1_down_t3_in  (r1_down_t3_in),
    .r1_up_t0_out   (r1_up_t0_out),
    .r1_up_t1_out   (r1_up_t1_out),
    .r1_up_t2_out   (r1_up_t2_out),
    .r1_up_t3_out   (r1_up_t3_out),
    .r1_down_t0_out (r1_down_t0_out),
    .r1_down_t1_out (r1_down_t1_out),
    .r1_down_t2_out (r1_down_t2_out),
    .r1_down_t3_out (r1_down_t3_out),
    .r2_up_t0_in    (r2_up_t0_in),
    .r2_up_t1_in    (r2_up_t1_in),
    .r2_up_t2_in    (r2_up_t2_in),
    .r2_up_t3_in    (r2_up_t3_in),
    .r2_down_t0_in  (r2_down_t0_in),
    .r2_down_t1_in  (r2_down_t1_in),
    .r2_down_t2_in  (r2_down_t2_in),
    .r2_down_t3_in  (r2_down_t3_in),
    .r2_up_t0_out   (r2_up_t0_out),
    .r2_up_t1_out   (r2_up_t1_out),
    .r2_up_t2_out   (r2_up_t2_out),
    .r2_up_t3_out   (r2_up_t3_out),
    .r2_down_t0_out (r2_down_t0_out),
    .r2_down_t1_out (r2_down_t1_out),
    .r2_down_t2_out (r2_down_t2_out),
    .r2_down_t3_out (r2_down_t3_out),
    .clk            (clk)
    );

  contol_switches contol_switches (
    .epsep         (epsep),
    .ep11          (ep11),
    .extended_pos  (extended_pos),
    .extended_neg  (extended_neg),
    .single_ep     (single_ep),
    .start         (start),
    .stop_neg      (stop_neg),
    .s2            (s2),
    .c22           (c22),
    .d18           (d[18]),
    .d35           (d[35]),
    .ep            (ep),
    .starter_neg   (starter_neg),
    .sep2          (sep2),
    .resume_btn    (resume_btn),
    .single_ep_btn (single_ep_btn),
    .start_btn     (start_btn),
    .stop_btn      (stop_btn),
    .extended_btn  (extended_btn)
    );

endmodule
