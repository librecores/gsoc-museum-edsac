module ccu_6
  (output reg ep,
   output reg ccu_ones,

   input wire ep0,
   input wire ep1,
   input wire ep2,
   input wire ep3,
   input wire ep4,
   input wire ep5,
   input wire ep6,
   input wire ep7,
   input wire ep8,
   input wire ep9,
   input wire ep10,
   input wire ep11,
   input wire ones1,
   input wire ones2,
   input wire ones4);

   // Body

endmodule // ccu_6
