module tank_dist_f2
  (output reg f2_down_f7_pos,
   output reg f2_up_f7_pos,
   output reg f2_down_f7_neg,
   output reg f2_up_f7_neg,
   output reg f2_down_f8_pos,
   output reg f2_up_f8_pos,
   output reg f2_down_f8_neg,
   output reg f2_up_f8_neg,
   output reg f2_down_t_in,
   output reg f2_up_t_in,
   output reg f2_down_t_out,
   output reg f2_up_t_out,

   input wire f2_down_dec_in,
   input wire f2_down_dec_out,
   input wire f2_up_dec_in,
   input wire f2_up_dec_out,
   input wire f7_pos,
   input wire f8_pos);

   // tank_dist to be instantiated here.
   
   // Body

endmodule // tank_dist_f2
