module main_ctrl
  (output reg ep_done,
   output reg g12,
   output reg g13,
   output reg r2,
   output reg s1,
   output reg s2,
   output reg sct_clear_gate,
   output reg sct_in_gate,
   output reg sct_one,

   input wire ep,
   input wire c17,
   input wire c21,
   input wire c26,
   input wire d0,
   input wire d18,
   input wire dv_d,
   input wire eng_mode_neg,
   input wire r_pulse,
   input wire single_ep,
   input wire stop_neg,
   input wire stop_one_a,
   input wire stop_one_b,
   input wire stop_one_c,
   input wire stop_one_d);

   // Body

endmodule // main_ctrl
