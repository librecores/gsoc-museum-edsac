module order_decoder2
  (output reg op1,
   output reg op2,
   output reg op3,
   output reg op4,
   output reg op5,
   output reg op6,
   output reg op7,
   output reg op8,

   input wire f13_pos,
   input wire f13_neg,
   input wire f14_pos,
   input wire f14_neg,
   input wire f15_pos,
   input wire f15_neg,
   input wire o_dy);

   // Body

endmodule // order_decoder2
