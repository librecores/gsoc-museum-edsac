module order_decoder2_3
  (output reg op_a,
   output reg op_b,
   output reg op_c,
   output reg op_delta,
   output reg op_g,
   output reg op_l,
   output reg op_v,
   output reg op_x,

   input wire f13_pos,
   input wire f13_neg,
   input wire f14_pos,
   input wire f14_neg,
   input wire f15_pos,
   input wire f15_neg,
   input wire o_dy_3);

   // One order_decoder2 to be instantiated.

endmodule // order_decoder2_3
