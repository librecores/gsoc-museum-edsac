module tank_dist
  (output reg rack_down_f7_pos,
   output reg rack_up_f7_pos,
   output reg rack_down_f7_neg,
   output reg rack_up_f7_neg,
   output reg rack_down_f8_pos,
   output reg rack_up_f8_pos,
   output reg rack_down_f8_neg,
   output reg rack_up_f8_neg,
   output reg rack_down_t_in,
   output reg rack_up_t_in,
   output reg rack_down_t_out,
   output reg rack_up_t_out,

   input wire rack_down_dec_in,
   input wire rack_down_dec_out,
   input wire rack_up_dec_in,
   input wire rack_up_dec_out,
   input wire f7_pos,
   input wire f8_pos);

   // Body

endmodule // tank_dist
