module order_decoder2_2
  (output reg op_blank,
   output reg op_d,
   output reg op_f,
   output reg op_h,
   output reg op_m,
   output reg op_n,
   output reg op_phi,
   output reg op_theta,

   input wire f13_pos,
   input wire f13_neg,
   input wire f14_pos,
   input wire f14_neg,
   input wire f15_pos,
   input wire f15_neg,
   input wire o_dy_2);

   // One order_decoder2 to be instantiated.

endmodule // order_decoder2_2
