module ccu_1
  (output reg odd_d35,
   output reg odd_d18,
   output reg odd_d0,
   output reg ev_d0,
   output reg ev_d1,
   output reg ev_d1_dz,
   output reg ev_d35,
   output reg g1_pos,
   output reg g1_neg,

   input wire d1,
   input wire d18,
   input wire d35,
   input wire da_n,
   input wire dy);

   // Body

endmodule // ccu_1
