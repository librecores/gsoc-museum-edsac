module tank_decoder1_f1
  (output reg f1_clk,
   output reg f1_down_dec_in,
   output reg f1_up_dec_in,
   output reg f1_down_dec_out,
   output reg f1_up_dec_out,
   output reg f1_down_t0_clr,
   output reg f1_up_t0_clr,
   output reg f1_down_t1_clr,
   output reg f1_up_t1_clr,
   output reg f1_down_t2_clr,
   output reg f1_up_t2_clr,
   output reg f1_down_t3_clr,
   output reg f1_up_t3_clr,
   output reg f1_mib,
   output reg f1_mob,

   input wire clk,
   input wire cls_neg,
   input wire f1_down_mob_t0,
   input wire f1_up_mob_t0,
   input wire f1_down_mob_t1,
   input wire f1_up_mob_t1,
   input wire f1_down_mob_t2,
   input wire f1_up_mob_t2,
   input wire f1_down_mob_t3,
   input wire f1_up_mob_t3,
   input wire f1_down_t0_in,
   input wire f1_up_t0_in,
   input wire f1_down_t1_in,
   input wire f1_up_t1_in,
   input wire f1_down_t2_in,
   input wire f1_up_t2_in,
   input wire f1_down_t3_in,
   input wire f1_up_t3_in,
   input wire f1_read,
   input wire f1_write,
   input wire f9_pos,
   input wire mib);

   // tank_decoder1 to be instantiated here.
   
   // Body

endmodule // tank_decoder1_f1
