module tank_decoder2_f2_down
  (output reg f2_down_t0_in,
   output reg f2_down_t0_out,
   output reg f2_down_t1_in,
   output reg f2_down_t1_out,
   output reg f2_down_t2_in,
   output reg f2_down_t2_out,
   output reg f2_down_t3_in,
   output reg f2_down_t3_out,

   input wire f2_down_f7_pos,
   input wire f2_down_f7_neg,
   input wire f2_down_f8_pos,
   input wire f2_down_f8_neg,
   input wire f2_down_t_in,
   input wire f2_down_t_out);

   // tank_decoder2 to be instantiated here.
   
   // Body

endmodule // tank_decoder2_f2_down
