module compl_collater(
                      // Outputs
                      adder_b,
                      // Inputs
                      clk, c2, c3, c4, c7, c9, ccu_ones, ev_d1_dz, g4_pos, g4_neg, mcand, mplier
                      );

   output reg adder_b;

   input wire clk;
   input wire c2;
   input wire c3;
   input wire c4;
   input wire c7;
   input wire c9;
   input wire ccu_ones;
   input wire ev_d1_dz;
   input wire g4_pos;
   input wire g4_neg;
   input wire multiplicand;
   input wire multiplier;

   // Body

endmodule // compl_collater
