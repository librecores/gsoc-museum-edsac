module order_coder
  (output reg c1,
   output reg c10,
   output reg c11,
   output reg c12,
   output reg c13,
   output reg c14,
   output reg c16,
   output reg c17,
   output reg c17a,
   output reg c18,
   output reg c19,
   output reg c2,
   output reg c20,
   output reg c21,
   output reg c22,
   output reg c24,
   output reg c25,
   output reg c26,
   output reg c27,
   output reg c3,
   output reg c4,
   output reg c5,
   output reg c6,
   output reg c7,
   output reg c8,
   output reg c9,

   input wire op_a,
   input wire op_b,
   input wire op_blank,
   input wire op_c,
   input wire op_d,
   input wire op_delta,
   input wire op_e,
   input wire op_erase,
   input wire op_f,
   input wire op_g,
   input wire op_h,
   input wire op_i,
   input wire op_j,
   input wire op_k,
   input wire op_l,
   input wire op_m,
   input wire op_n,
   input wire op_o,
   input wire op_p,
   input wire op_phi,
   input wire op_pi,
   input wire op_q,
   input wire op_r,
   input wire op_s,
   input wire op_t,
   input wire op_theta,
   input wire op_u,
   input wire op_v,
   input wire op_w,
   input wire op_x,
   input wire op_y,
   input wire op_z,
   input wire starter,
   input wire starter_neg,
   input wire extended_neg);

   // Body

endmodule // order_coder
