module memory_f2_down_0
  (output reg monitor13,
   output reg f2_down_mob_t0,

   input wire f2_clk,
   input wire f2_mib,
   input wire f2_down_t0_clr,
   input wire f2_down_t0_in,
   input wire f2_down_t0_out);

   // Atomic dleay_line module to be instantiated here 
   // with 1.152ms delay for circulation of 16 full 
   // words or 32 short words (instructions).

   // Body

endmodule // memory_f2_down_0
