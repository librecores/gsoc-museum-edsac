module sequence_ctrl_tank
  (output reg sct,

   input wire clk,
   input wire g12,
   input wire sct_clear_gate,
   input wire sct_in_gate,
   input wire sct_one,
   input wire ungated_order,
   input wire reset_sct);

   // One half adder to be instantiated 
   // along with half cycle delay.

   // Body

endmodule // sequence_ctrl_tank
