module memory_r1_up_0
  (output reg monitor17,
   output reg r1_up_mob_t0,

   input wire r1_clk,
   input wire r1_mib,
   input wire r1_up_t0_clr,
   input wire r1_up_t0_in,
   input wire r1_up_t0_out);

   // Atomic dleay_line module to be instantiated here 
   // with 1.152ms delay for circulation of 16 full 
   // words or 32 short words (instructions).

   // Body

endmodule // memory_r1_up_0
