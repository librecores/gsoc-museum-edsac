/* Module for Control Switches Unit.
 */

module contol_switches (
  output wire epsep,
  output wire ep11,
  output wire extended_pos,
  output wire extended_neg,
  output wire single_ep,
  output wire start,
  output wire stop_neg,

  input wire  s2,
  input wire  c22,
  input wire  d18,
  input wire  d35,
  input wire  ep,
  input wire  starter_neg,
  input wire  sep2
  );

endmodule
