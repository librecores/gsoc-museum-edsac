/* Top Level L0 EDSAC module.
 */

module edsac (
  input wire clk
  );

  wire        f1_down_mob_t0;
  wire        f1_up_mob_t0;
  wire        f1_down_mob_t1;
  wire        f1_up_mob_t1;
  wire        f1_down_mob_t2;
  wire        f1_up_mob_t2;
  wire        f1_down_mob_t3;
  wire        f1_up_mob_t3;
  wire        f2_down_mob_t0;
  wire        f2_up_mob_t0;
  wire        f2_down_mob_t1;
  wire        f2_up_mob_t1;
  wire        f2_down_mob_t2;
  wire        f2_up_mob_t2;
  wire        f2_down_mob_t3;
  wire        f2_up_mob_t3;
  wire        r1_down_mob_t0;
  wire        r1_up_mob_t0;
  wire        r1_down_mob_t1;
  wire        r1_up_mob_t1;
  wire        r1_down_mob_t2;
  wire        r1_up_mob_t2;
  wire        r1_down_mob_t3;
  wire        r1_up_mob_t3;
  wire        r2_down_mob_t0;
  wire        r2_up_mob_t0;
  wire        r2_down_mob_t1;
  wire        r2_up_mob_t1;
  wire        r2_down_mob_t2;
  wire        r2_up_mob_t2;
  wire        r2_down_mob_t3;
  wire        r2_up_mob_t3;
  wire        f1_mib;
  wire        f2_mib;
  wire        r1_mib;
  wire        r2_mib;
  wire        f1_down_t0_clr;
  wire        f1_up_t0_clr;
  wire        f1_down_t1_clr;
  wire        f1_up_t1_clr;
  wire        f1_down_t2_clr;
  wire        f1_up_t2_clr;
  wire        f1_down_t3_clr;
  wire        f1_up_t3_clr;
  wire        f2_down_t0_clr;
  wire        f2_up_t0_clr;
  wire        f2_down_t1_clr;
  wire        f2_up_t1_clr;
  wire        f2_down_t2_clr;
  wire        f2_up_t2_clr;
  wire        f2_down_t3_clr;
  wire        f2_up_t3_clr;
  wire        r1_down_t0_clr;
  wire        r1_up_t0_clr;
  wire        r1_down_t1_clr;
  wire        r1_up_t1_clr;
  wire        r1_down_t2_clr;
  wire        r1_up_t2_clr;
  wire        r1_down_t3_clr;
  wire        r1_up_t3_clr;
  wire        r2_down_t0_clr;
  wire        r2_up_t0_clr;
  wire        r2_down_t1_clr;
  wire        r2_up_t1_clr;
  wire        r2_down_t2_clr;
  wire        r2_up_t2_clr;
  wire        r2_down_t3_clr;
  wire        r2_up_t3_clr;
  wire        f1_up_t0_in;
  wire        f1_up_t1_in;
  wire        f1_up_t2_in;
  wire        f1_up_t3_in;
  wire        f1_down_t0_in;
  wire        f1_down_t1_in;
  wire        f1_down_t2_in;
  wire        f1_down_t3_in;
  wire        f1_up_t0_out;
  wire        f1_up_t1_out;
  wire        f1_up_t2_out;
  wire        f1_up_t3_out;
  wire        f1_down_t0_out;
  wire        f1_down_t1_out;
  wire        f1_down_t2_out;
  wire        f1_down_t3_out;
  wire        f2_up_t0_in;
  wire        f2_up_t1_in;
  wire        f2_up_t2_in;
  wire        f2_up_t3_in;
  wire        f2_down_t0_in;
  wire        f2_down_t1_in;
  wire        f2_down_t2_in;
  wire        f2_down_t3_in;
  wire        f2_up_t0_out;
  wire        f2_up_t1_out;
  wire        f2_up_t2_out;
  wire        f2_up_t3_out;
  wire        f2_down_t0_out;
  wire        f2_down_t1_out;
  wire        f2_down_t2_out;
  wire        f2_down_t3_out;
  wire        r1_up_t0_in;
  wire        r1_up_t1_in;
  wire        r1_up_t2_in;
  wire        r1_up_t3_in;
  wire        r1_down_t0_in;
  wire        r1_down_t1_in;
  wire        r1_down_t2_in;
  wire        r1_down_t3_in;
  wire        r1_up_t0_out;
  wire        r1_up_t1_out;
  wire        r1_up_t2_out;
  wire        r1_up_t3_out;
  wire        r1_down_t0_out;
  wire        r1_down_t1_out;
  wire        r1_down_t2_out;
  wire        r1_down_t3_out;
  wire        r2_up_t0_in;
  wire        r2_up_t1_in;
  wire        r2_up_t2_in;
  wire        r2_up_t3_in;
  wire        r2_down_t0_in;
  wire        r2_down_t1_in;
  wire        r2_down_t2_in;
  wire        r2_down_t3_in;
  wire        r2_up_t0_out;
  wire        r2_up_t1_out;
  wire        r2_up_t2_out;
  wire        r2_up_t3_out;
  wire        r2_down_t0_out;
  wire        r2_down_t1_out;
  wire        r2_down_t2_out;
  wire        r2_down_t3_out;
  wire [35:0] d;

  digit_pulse_generator digit_pulse_generator (
    .digit_pulse (d[35:0]),
    
    .clk (clk)
    );

  memory_top memory_top (
    // TODO: monitors are for displaying Tank contents and are not connected for now.
    .monitor1       (),
    .monitor2       (),
    .monitor3       (),
    .monitor4       (),
    .monitor5       (),
    .monitor6       (),
    .monitor7       (),
    .monitor8       (),
    .monitor9       (),
    .monitor10      (),
    .monitor11      (),
    .monitor12      (),
    .monitor13      (),
    .monitor14      (),
    .monitor15      (),
    .monitor16      (),
    .monitor17      (),
    .monitor18      (),
    .monitor19      (),
    .monitor20      (),
    .monitor21      (),
    .monitor22      (),
    .monitor23      (),
    .monitor24      (),
    .monitor25      (),
    .monitor26      (),
    .monitor27      (),
    .monitor28      (),
    .monitor29      (),
    .monitor30      (),
    .monitor31      (),
    .monitor32      (),
    .f1_down_mob_t0 (f1_down_mob_t0),
    .f1_up_mob_t0   (f1_up_mob_t0),
    .f1_down_mob_t1 (f1_down_mob_t1),
    .f1_up_mob_t1   (f1_up_mob_t1),
    .f1_down_mob_t2 (f1_down_mob_t2),
    .f1_up_mob_t2   (f1_up_mob_t2),
    .f1_down_mob_t3 (f1_down_mob_t3),
    .f1_up_mob_t3   (f1_up_mob_t3),
    .f2_down_mob_t0 (f2_down_mob_t0),
    .f2_up_mob_t0   (f2_up_mob_t0),
    .f2_down_mob_t1 (f2_down_mob_t1),
    .f2_up_mob_t1   (f2_up_mob_t1),
    .f2_down_mob_t2 (f2_down_mob_t2),
    .f2_up_mob_t2   (f2_up_mob_t2),
    .f2_down_mob_t3 (f2_down_mob_t3),
    .f2_up_mob_t3   (f2_up_mob_t3),
    .r1_down_mob_t0 (r1_down_mob_t0),
    .r1_up_mob_t0   (r1_up_mob_t0),
    .r1_down_mob_t1 (r1_down_mob_t1),
    .r1_up_mob_t1   (r1_up_mob_t1),
    .r1_down_mob_t2 (r1_down_mob_t2),
    .r1_up_mob_t2   (r1_up_mob_t2),
    .r1_down_mob_t3 (r1_down_mob_t3),
    .r1_up_mob_t3   (r1_up_mob_t3),
    .r2_down_mob_t0 (r2_down_mob_t0),
    .r2_up_mob_t0   (r2_up_mob_t0),
    .r2_down_mob_t1 (r2_down_mob_t1),
    .r2_up_mob_t1   (r2_up_mob_t1),
    .r2_down_mob_t2 (r2_down_mob_t2),
    .r2_up_mob_t2   (r2_up_mob_t2),
    .r2_down_mob_t3 (r2_down_mob_t3),
    .r2_up_mob_t3   (r2_up_mob_t3),

    .f1_mib         (f1_mib),
    .f2_mib         (f2_mib),
    .r1_mib         (r1_mib),
    .r2_mib         (r2_mib),
    .f1_down_t0_clr (f1_down_t0_clr),
    .f1_up_t0_clr   (f1_up_t0_clr),
    .f1_down_t1_clr (f1_down_t1_clr),
    .f1_up_t1_clr   (f1_up_t1_clr),
    .f1_down_t2_clr (f1_down_t2_clr),
    .f1_up_t2_clr   (f1_up_t2_clr),
    .f1_down_t3_clr (f1_down_t3_clr),
    .f1_up_t3_clr   (f1_up_t3_clr),
    .f2_down_t0_clr (f2_down_t0_clr),
    .f2_up_t0_clr   (f2_up_t0_clr),
    .f2_down_t1_clr (f2_down_t1_clr),
    .f2_up_t1_clr   (f2_up_t1_clr),
    .f2_down_t2_clr (f2_down_t2_clr),
    .f2_up_t2_clr   (f2_up_t2_clr),
    .f2_down_t3_clr (f2_down_t3_clr),
    .f2_up_t3_clr   (f2_up_t3_clr),
    .r1_down_t0_clr (r1_down_t0_clr),
    .r1_up_t0_clr   (r1_up_t0_clr),
    .r1_down_t1_clr (r1_down_t1_clr),
    .r1_up_t1_clr   (r1_up_t1_clr),
    .r1_down_t2_clr (r1_down_t2_clr),
    .r1_up_t2_clr   (r1_up_t2_clr),
    .r1_down_t3_clr (r1_down_t3_clr),
    .r1_up_t3_clr   (r1_up_t3_clr),
    .r2_down_t0_clr (r2_down_t0_clr),
    .r2_up_t0_clr   (r2_up_t0_clr),
    .r2_down_t1_clr (r2_down_t1_clr),
    .r2_up_t1_clr   (r2_up_t1_clr),
    .r2_down_t2_clr (r2_down_t2_clr),
    .r2_up_t2_clr   (r2_up_t2_clr),
    .r2_down_t3_clr (r2_down_t3_clr),
    .r2_up_t3_clr   (r2_up_t3_clr),
    .f1_up_t0_in    (f1_up_t0_in),
    .f1_up_t1_in    (f1_up_t1_in),
    .f1_up_t2_in    (f1_up_t2_in),
    .f1_up_t3_in    (f1_up_t3_in),
    .f1_down_t0_in  (f1_down_t0_in),
    .f1_down_t1_in  (f1_down_t1_in),
    .f1_down_t2_in  (f1_down_t2_in),
    .f1_down_t3_in  (f1_down_t3_in),
    .f1_up_t0_out   (f1_up_t0_out),
    .f1_up_t1_out   (f1_up_t1_out),
    .f1_up_t2_out   (f1_up_t2_out),
    .f1_up_t3_out   (f1_up_t3_out),
    .f1_down_t0_out (f1_down_t0_out),
    .f1_down_t1_out (f1_down_t1_out),
    .f1_down_t2_out (f1_down_t2_out),
    .f1_down_t3_out (f1_down_t3_out),
    .f2_up_t0_in    (f2_up_t0_in),
    .f2_up_t1_in    (f2_up_t1_in),
    .f2_up_t2_in    (f2_up_t2_in),
    .f2_up_t3_in    (f2_up_t3_in),
    .f2_down_t0_in  (f2_down_t0_in),
    .f2_down_t1_in  (f2_down_t1_in),
    .f2_down_t2_in  (f2_down_t2_in),
    .f2_down_t3_in  (f2_down_t3_in),
    .f2_up_t0_out   (f2_up_t0_out),
    .f2_up_t1_out   (f2_up_t1_out),
    .f2_up_t2_out   (f2_up_t2_out),
    .f2_up_t3_out   (f2_up_t3_out),
    .f2_down_t0_out (f2_down_t0_out),
    .f2_down_t1_out (f2_down_t1_out),
    .f2_down_t2_out (f2_down_t2_out),
    .f2_down_t3_out (f2_down_t3_out),
    .r1_up_t0_in    (r1_up_t0_in),
    .r1_up_t1_in    (r1_up_t1_in),
    .r1_up_t2_in    (r1_up_t2_in),
    .r1_up_t3_in    (r1_up_t3_in),
    .r1_down_t0_in  (r1_down_t0_in),
    .r1_down_t1_in  (r1_down_t1_in),
    .r1_down_t2_in  (r1_down_t2_in),
    .r1_down_t3_in  (r1_down_t3_in),
    .r1_up_t0_out   (r1_up_t0_out),
    .r1_up_t1_out   (r1_up_t1_out),
    .r1_up_t2_out   (r1_up_t2_out),
    .r1_up_t3_out   (r1_up_t3_out),
    .r1_down_t0_out (r1_down_t0_out),
    .r1_down_t1_out (r1_down_t1_out),
    .r1_down_t2_out (r1_down_t2_out),
    .r1_down_t3_out (r1_down_t3_out),
    .r2_up_t0_in    (r2_up_t0_in),
    .r2_up_t1_in    (r2_up_t1_in),
    .r2_up_t2_in    (r2_up_t2_in),
    .r2_up_t3_in    (r2_up_t3_in),
    .r2_down_t0_in  (r2_down_t0_in),
    .r2_down_t1_in  (r2_down_t1_in),
    .r2_down_t2_in  (r2_down_t2_in),
    .r2_down_t3_in  (r2_down_t3_in),
    .r2_up_t0_out   (r2_up_t0_out),
    .r2_up_t1_out   (r2_up_t1_out),
    .r2_up_t2_out   (r2_up_t2_out),
    .r2_up_t3_out   (r2_up_t3_out),
    .r2_down_t0_out (r2_down_t0_out),
    .r2_down_t1_out (r2_down_t1_out),
    .r2_down_t2_out (r2_down_t2_out),
    .r2_down_t3_out (r2_down_t3_out),
    .clk            (clk)
    );

endmodule
