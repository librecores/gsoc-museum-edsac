module half_adder(
                  // Outputs
                  sum, carry,
                  // Inputs
                  clk, operand_a, operand_b
                  );

   output reg sum;
   output reg carry;

   input wire clk;
   input wire operand_a;
   input wire operand_b;

   // Body

endmodule // half_adder
