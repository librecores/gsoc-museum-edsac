module tank_decoder1_r1
  (output reg r1_clk,
   output reg r1_down_dec_in,
   output reg r1_up_dec_in,
   output reg r1_down_dec_out,
   output reg r1_up_dec_out,
   output reg r1_down_t0_clr,
   output reg r1_up_t0_clr,
   output reg r1_down_t1_clr,
   output reg r1_up_t1_clr,
   output reg r1_down_t2_clr,
   output reg r1_up_t2_clr,
   output reg r1_down_t3_clr,
   output reg r1_up_t3_clr,
   output reg r1_mib,
   output reg r1_mob,

   input wire clk,
   input wire cls_neg,
   input wire r1_down_mob_t0,
   input wire r1_up_mob_t0,
   input wire r1_down_mob_t1,
   input wire r1_up_mob_t1,
   input wire r1_down_mob_t2,
   input wire r1_up_mob_t2,
   input wire r1_down_mob_t3,
   input wire r1_up_mob_t3,
   input wire r1_down_t0_in,
   input wire r1_up_t0_in,
   input wire r1_down_t1_in,
   input wire r1_up_t1_in,
   input wire r1_down_t2_in,
   input wire r1_up_t2_in,
   input wire r1_down_t3_in,
   input wire r1_up_t3_in,
   input wire r1_read,
   input wire r1_write,
   input wire f9_pos,
   input wire mib);

   // tank_decoder1 to be instantiated here.
   
   // Body

endmodule // tank_decoder1_r1
