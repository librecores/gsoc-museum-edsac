module adder(
             // Outputs
             adder_sum,
             // Inputs
             clk, adder_a, adder_b, ev_d1
             );

   output adder_sum;

   input wire clk;
   input wire adder_a;
   input wire adder_b;
   input wire ev_d1;

   // Two half adders to be instantiated here -
   // one with feedback and the other without.

   // Body
   
endmodule // adder
