module tank_flash
  (output reg f1_pos,
   output reg f1_neg,
   output reg f10_pos,
   output reg f11_pos,
   output reg f2_pos,
   output reg f7_pos,
   output reg f8_pos,
   output reg f9_pos,

   input wire d19,
   input wire d20,
   input wire d25,
   input wire d26,
   input wire d27,
   input wire d28,
   input wire d29,
   input wire epsep,
   input wire g12,
   input wire order_sct);

   // Body

endmodule // tank_flash
