module tank_decoder1_f2
  (output reg f2_clk,
   output reg f2_down_dec_in,
   output reg f2_up_dec_in,
   output reg f2_down_dec_out,
   output reg f2_up_dec_out,
   output reg f2_down_t0_clr,
   output reg f2_up_t0_clr,
   output reg f2_down_t1_clr,
   output reg f2_up_t1_clr,
   output reg f2_down_t2_clr,
   output reg f2_up_t2_clr,
   output reg f2_down_t3_clr,
   output reg f2_up_t3_clr,
   output reg f2_mib,
   output reg f2_mob,

   input wire clk,
   input wire cls_neg,
   input wire f2_down_mob_t0,
   input wire f2_up_mob_t0,
   input wire f2_down_mob_t1,
   input wire f2_up_mob_t1,
   input wire f2_down_mob_t2,
   input wire f2_up_mob_t2,
   input wire f2_down_mob_t3,
   input wire f2_up_mob_t3,
   input wire f2_down_t0_in,
   input wire f2_up_t0_in,
   input wire f2_down_t1_in,
   input wire f2_up_t1_in,
   input wire f2_down_t2_in,
   input wire f2_up_t2_in,
   input wire f2_down_t3_in,
   input wire f2_up_t3_in,
   input wire f2_read,
   input wire f2_write,
   input wire f9_pos,
   input wire mib);

   // tank_decoder1 to be instantiated here.
   
   // Body

endmodule // tank_decoder1_f2
