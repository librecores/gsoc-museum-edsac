module tank_decoder2
  (output reg rack_loc_t0_in,
   output reg rack_loc_t0_out,
   output reg rack_loc_t1_in,
   output reg rack_loc_t1_out,
   output reg rack_loc_t2_in,
   output reg rack_loc_t2_out,
   output reg rack_loc_t3_in,
   output reg rack_loc_t3_out,

   input wire rack_loc_f7_pos,
   input wire rack_loc_f7_neg,
   input wire rack_loc_f8_pos,
   input wire rack_loc_f8_neg,
   input wire rack_loc_t_in,
   input wire rack_loc_t_out);

   // Body

endmodule // tank_decoder2
