module ccu_2
  (output reg zero_d0,
   output reg da_m,
   output reg ds,
   output reg g8,

   input wire c5,
   input wire c6,
   input wire c7,
   input wire d35,
   input wire da,
   input wire ev_d0,
   input wire mcand_in,
   input wire s2);

   // Body

endmodule // ccu_2
