module multiplicand(
                    // Outputs
                    da_n, mcand, mcand_in,
                    // Inputs
                    clk, c1, c21, da_m, g11_neg, g12, g13, g2_pos, g2_neg, g3_pos, g6_pos, mib
                    );

   output reg da_n;
   output reg mcand;
   output reg mcand_in;

   input wire clk;
   input wire c1;
   input wire c21;
   input wire da_m;
   input wire g11_neg;
   input wire g12;
   input wire g13;
   input wire g2_pos;
   input wire g2_neg;
   input wire g3_pos;
   input wire g6_pos;
   input wire mib;

   // Body

endmodule // multiplicand
