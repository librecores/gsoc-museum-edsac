module ccu_9_11
  (output reg ep6,
   output reg ep7,
   output reg g9_neg,
   output reg g10_neg,
   output reg g11_neg,

   input wire c18,
   input wire c19,
   input wire c20,
   input wire ev_d0,
   input wire odd_d0,
   input wire r2,
   input wire s2,
   input wire op_u);

   // Body

endmodule // ccu_9_11
