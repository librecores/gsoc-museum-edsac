module acc_shift_i(
                   // Outputs
                   mob8, x1, x2, x3, x4,
                   // Inputs
                   clk, acc, c19, c7, c8, d17, d35, f1_neg, g5
                   );

   output reg mob8;
   output reg x1;
   output reg x2;
   output reg x3;
   output reg x4;

   input wire clk;
   input wire acc;
   input wire c19;
   input wire c7;
   input wire c8;
   input wire d17;
   input wire d35;
   input wire f1_neg;
   input wire g5;

   // Body

endmodule // acc_shift_i
