module compl_collater
  (output reg adder_b,

   input wire clk,
   input wire c2,
   input wire c3,
   input wire c4,
   input wire c7,
   input wire c9,
   input wire ccu_ones,
   input wire ev_d1_dz,
   input wire g4_pos,
   input wire g4_neg,
   input wire mcand,
   input wire mplier);

   // Body

endmodule // compl_collater
