module ccu_5
  (output reg ep0,
   output reg ones4,

   input wire c9,
   input wire c12,
   input wire c13,
   input wire d18,
   input wire ep_done,
   input wire ev_d0,
   input wire extended_neg,
   input wire odd_d0,
   input wire s2);

   // Body

endmodule // ccu_5
