/* Top module for Memory L1 subsystem.
 */

module memory_top (
  output wire [575:0] monitor1,
  output wire [575:0] monitor2,
  output wire [575:0] monitor3,
  output wire [575:0] monitor4,
  output wire [575:0] monitor5,
  output wire [575:0] monitor6,
  output wire [575:0] monitor7,
  output wire [575:0] monitor8,
  output wire [575:0] monitor9,
  output wire [575:0] monitor10,
  output wire [575:0] monitor11,
  output wire [575:0] monitor12,
  output wire [575:0] monitor13,
  output wire [575:0] monitor14,
  output wire [575:0] monitor15,
  output wire [575:0] monitor16,
  output wire [575:0] monitor17,
  output wire [575:0] monitor18,
  output wire [575:0] monitor19,
  output wire [575:0] monitor20,
  output wire [575:0] monitor21,
  output wire [575:0] monitor22,
  output wire [575:0] monitor23,
  output wire [575:0] monitor24,
  output wire [575:0] monitor25,
  output wire [575:0] monitor26,
  output wire [575:0] monitor27,
  output wire [575:0] monitor28,
  output wire [575:0] monitor29,
  output wire [575:0] monitor30,
  output wire [575:0] monitor31,
  output wire [575:0] monitor32,
  output wire f1_down_mob_t0,
  output wire f1_up_mob_t0,
  output wire f1_down_mob_t1,
  output wire f1_up_mob_t1,
  output wire f1_down_mob_t2,
  output wire f1_up_mob_t2,
  output wire f1_down_mob_t3,
  output wire f1_up_mob_t3,
  output wire f2_down_mob_t0,
  output wire f2_up_mob_t0,
  output wire f2_down_mob_t1,
  output wire f2_up_mob_t1,
  output wire f2_down_mob_t2,
  output wire f2_up_mob_t2,
  output wire f2_down_mob_t3,
  output wire f2_up_mob_t3,
  output wire r1_down_mob_t0,
  output wire r1_up_mob_t0,
  output wire r1_down_mob_t1,
  output wire r1_up_mob_t1,
  output wire r1_down_mob_t2,
  output wire r1_up_mob_t2,
  output wire r1_down_mob_t3,
  output wire r1_up_mob_t3,
  output wire r2_down_mob_t0,
  output wire r2_up_mob_t0,
  output wire r2_down_mob_t1,
  output wire r2_up_mob_t1,
  output wire r2_down_mob_t2,
  output wire r2_up_mob_t2,
  output wire r2_down_mob_t3,
  output wire r2_up_mob_t3,

  input wire  f1_mib,
  input wire  f2_mib,
  input wire  r1_mib,
  input wire  r2_mib,
  input wire  f1_down_t0_clr,
  input wire  f1_up_t0_clr,
  input wire  f1_down_t1_clr,
  input wire  f1_up_t1_clr,
  input wire  f1_down_t2_clr,
  input wire  f1_up_t2_clr,
  input wire  f1_down_t3_clr,
  input wire  f1_up_t3_clr,
  input wire  f2_down_t0_clr,
  input wire  f2_up_t0_clr,
  input wire  f2_down_t1_clr,
  input wire  f2_up_t1_clr,
  input wire  f2_down_t2_clr,
  input wire  f2_up_t2_clr,
  input wire  f2_down_t3_clr,
  input wire  f2_up_t3_clr,
  input wire  r1_down_t0_clr,
  input wire  r1_up_t0_clr,
  input wire  r1_down_t1_clr,
  input wire  r1_up_t1_clr,
  input wire  r1_down_t2_clr,
  input wire  r1_up_t2_clr,
  input wire  r1_down_t3_clr,
  input wire  r1_up_t3_clr,
  input wire  r2_down_t0_clr,
  input wire  r2_up_t0_clr,
  input wire  r2_down_t1_clr,
  input wire  r2_up_t1_clr,
  input wire  r2_down_t2_clr,
  input wire  r2_up_t2_clr,
  input wire  r2_down_t3_clr,
  input wire  r2_up_t3_clr,
  input wire  f1_up_t0_in,
  input wire  f1_up_t1_in,
  input wire  f1_up_t2_in,
  input wire  f1_up_t3_in,
  input wire  f1_down_t0_in,
  input wire  f1_down_t1_in,
  input wire  f1_down_t2_in,
  input wire  f1_down_t3_in,
  input wire  f1_up_t0_out,
  input wire  f1_up_t1_out,
  input wire  f1_up_t2_out,
  input wire  f1_up_t3_out,
  input wire  f1_down_t0_out,
  input wire  f1_down_t1_out,
  input wire  f1_down_t2_out,
  input wire  f1_down_t3_out,
  input wire  f2_up_t0_in,
  input wire  f2_up_t1_in,
  input wire  f2_up_t2_in,
  input wire  f2_up_t3_in,
  input wire  f2_down_t0_in,
  input wire  f2_down_t1_in,
  input wire  f2_down_t2_in,
  input wire  f2_down_t3_in,
  input wire  f2_up_t0_out,
  input wire  f2_up_t1_out,
  input wire  f2_up_t2_out,
  input wire  f2_up_t3_out,
  input wire  f2_down_t0_out,
  input wire  f2_down_t1_out,
  input wire  f2_down_t2_out,
  input wire  f2_down_t3_out,
  input wire  r1_up_t0_in,
  input wire  r1_up_t1_in,
  input wire  r1_up_t2_in,
  input wire  r1_up_t3_in,
  input wire  r1_down_t0_in,
  input wire  r1_down_t1_in,
  input wire  r1_down_t2_in,
  input wire  r1_down_t3_in,
  input wire  r1_up_t0_out,
  input wire  r1_up_t1_out,
  input wire  r1_up_t2_out,
  input wire  r1_up_t3_out,
  input wire  r1_down_t0_out,
  input wire  r1_down_t1_out,
  input wire  r1_down_t2_out,
  input wire  r1_down_t3_out,
  input wire  r2_up_t0_in,
  input wire  r2_up_t1_in,
  input wire  r2_up_t2_in,
  input wire  r2_up_t3_in,
  input wire  r2_down_t0_in,
  input wire  r2_down_t1_in,
  input wire  r2_down_t2_in,
  input wire  r2_down_t3_in,
  input wire  r2_up_t0_out,
  input wire  r2_up_t1_out,
  input wire  r2_up_t2_out,
  input wire  r2_up_t3_out,
  input wire  r2_down_t0_out,
  input wire  r2_down_t1_out,
  input wire  r2_down_t2_out,
  input wire  r2_down_t3_out,
  input wire  clk
  );

endmodule
