module tank_decoder2_r1_down
  (output reg r1_down_t0_in,
   output reg r1_down_t0_out,
   output reg r1_down_t1_in,
   output reg r1_down_t1_out,
   output reg r1_down_t2_in,
   output reg r1_down_t2_out,
   output reg r1_down_t3_in,
   output reg r1_down_t3_out,

   input wire r1_down_f7_pos,
   input wire r1_down_f7_neg,
   input wire r1_down_f8_pos,
   input wire r1_down_f8_neg,
   input wire r1_down_t_in,
   input wire r1_down_t_out);

   // tank_decoder2 to be instantiated here.
   
   // Body

endmodule // tank_decoder2_r1_down
