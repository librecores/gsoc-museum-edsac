module delay_line
  (output reg data_out,

   input wire clk,
   input wire data_in);

   // Body

endmodule // delay_line
