module adder
  (output reg adder_sum,

   input wire clk,
   input wire adder_a,
   input wire adder_b,
   input wire ev_d1);

   // Two half adders to be instantiated here - 
   // one with feedback and other without.
   
   // Body

endmodule // adder
