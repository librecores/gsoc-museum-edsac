module transfer
  (output reg mib,
   output reg mob,

   input wire clk,
   input wire f1_pos,
   input wire f1_mob,
   input wire f2_pos,
   input wire f2_mob,
   input wire mob8,
   input wire mob9,
   input wire mob10,
   input wire mob11,
   input wire r1_mob,
   input wire r2_mob);

   // Body

endmodule // transfer
