module tank_decoder2_f1_up
  (output reg f1_up_t0_in,
   output reg f1_up_t0_out,
   output reg f1_up_t1_in,
   output reg f1_up_t1_out,
   output reg f1_up_t2_in,
   output reg f1_up_t2_out,
   output reg f1_up_t3_in,
   output reg f1_up_t3_out,

   input wire f1_up_f7_pos,
   input wire f1_up_f7_neg,
   input wire f1_up_f8_pos,
   input wire f1_up_f8_neg,
   input wire f1_up_t_in,
   input wire f1_up_t_out);

   // tank_decoder2 to be instantiated here.
   
   // Body

endmodule // tank_decoder2_f1_up
