module ccu_10
  (output reg dv,
   output reg ep5,
   output reg jump_uc,
   output reg stop_one_b,

   input wire c10,
   input wire c25,
   input wire d35,
   input wire dv_d,
   input wire ep_done,
   input wire ev_d0,
   input wire extended_pos,
   input wire odd_d0,
   input wire op_j,
   input wire s2);

   // Body

endmodule // ccu_10
