module order_flash
  (output reg f13_pos,
   output reg f13_neg,
   output reg f14_pos,
   output reg f14_neg,
   output reg f15_pos,
   output reg f15_neg,
   output reg f16_pos,
   output reg f16_neg,
   output reg f17_pos,
   output reg f17_neg,
   output reg order_flash_rdy,

   input wire d31,
   input wire d32,
   input wire d33,
   input wire d34,
   input wire d35,
   input wire epsep,
   input wire order);

   // Body

endmodule // order_flash
