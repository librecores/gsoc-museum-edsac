module tank_decoder0
  (output reg f1_read,
   output reg f1_write,
   output reg f2_read,
   output reg f2_write,
   output reg r1_read,
   output reg r1_write,
   output reg r2_read,
   output reg r2_write,

   input wire c17a,
   input wire f10_pos,
   input wire f11_pos,
   input wire cu_gate_pos);

   // Body

endmodule // tank_decoder0
