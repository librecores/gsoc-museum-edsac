module multiplicand
  (output reg da_n,
   output reg mcand,
   output reg mcand_in,

   input wire clk,
   input wire c1,
   input wire c21,
   input wire da_m,
   input wire g11_neg,
   input wire g12,
   input wire g13,
   input wire g2_pos,
   input wire g2_neg,
   input wire g3_pos,
   input wire g6_pos,
   input wire mib);

   // Body

endmodule // multiplicand
