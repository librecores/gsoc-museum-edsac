module order_decoder1
  (output reg o_dy_0,
   output reg o_dy_1,
   output reg o_dy_2,
   output reg o_dy_3,

   input wire f16_pos,
   input wire f16_neg,
   input wire f17_pos,
   input wire f17_neg,
   input wire order_flash_rdy);

   // Body

endmodule // order_decoder1
