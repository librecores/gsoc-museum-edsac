module timing_ctrl_shift
  (output reg seventy_d35,
   output reg da,
   output reg dx,
   output reg dy,
   output reg g2_pos,
   output reg g2_neg,

   input wire clk,
   input wire c5,
   input wire c6,
   input wire zero_d0,
   input wire d35);

   // Body

endmodule // timing_ctrl_shift
