module multiplier
  (output reg dx_m,
   output reg ep4,
   output reg mpier,

   input wire clk,
   input wire c18,
   input wire d35,
   input wire dx,
   input wire g10_neg,
   input wire mib,
   input wire r2);

   // Body

endmodule // multiplier

