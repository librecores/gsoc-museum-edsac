module memory_f2_up_3
  (output reg monitor12,
   output reg f2_up_mob_t3,

   input wire f2_clk,
   input wire f2_mib,
   input wire f2_up_t3_clr,
   input wire f2_up_t3_in,
   input wire f2_up_t3_out);

   // Atomic dleay_line module to be instantiated here 
   // with 1.152ms delay for circulation of 16 full 
   // words or 32 short words (instructions).

   // Body

endmodule // memory_f2_up_3
