module order_decoder2_0
  (output reg op_e,
   output reg op_p,
   output reg op_q,
   output reg op_r,
   output reg op_t,
   output reg op_u,
   output reg op_w,
   output reg op_y,

   input wire f13_pos,
   input wire f13_neg,
   input wire f14_pos,
   input wire f14_neg,
   input wire f15_pos,
   input wire f15_neg,
   input wire o_dy_0);

   // One order_decoder2 to be instantiated.

endmodule // order_decoder2_0
