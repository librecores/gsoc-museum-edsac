module multiplier(
                  // Outputs
                  dx_m, ep4, mpier,
                  // Inputs
                  clk, c18, d35, dx, g10_neg, mib, r2
                  );

   output reg dx_m;
   output reg ep4;
   output reg mpier;

   input wire clk;
   input wire c18;
   input wire d35;
   input wire dx;
   input wire g10_neg;
   input wire mib;
   input wire r2;

   // Body

endmodule // multiplier
